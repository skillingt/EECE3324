/*
 * Taylor Skilling
 * Will Johnson
 * 12/14/2016
 * EECE 3324
 *
 * mux3to1.v -- 32-bit 3:1 mux for X stage 
 */

module mux3to1(I0, I1, I2, S0, A);
input [31:0] I0, I1, I2; 
input [1:0] S0;          
output reg [31:0] A;    

initial
begin
    A = 0;
end
  
always @ (I0 or I1 or I2 or S0) begin
    case(S0)
      2'b00: begin
        A <= I0;
      end
      2'b01: begin
        A <= I1;
      end
      2'b10: begin
        A <= I2;
      end
    endcase
  end

endmodule
